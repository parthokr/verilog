module addOne (
    input wire [6:0] I,
    output wire [6:0] O
);
    assign O = I + 1'b1;
endmodule